module circuit_a(
    // Declare inputs
    // Declare Y output
);

    // Enter logic equation here
    (C | D) & (~C | D) & (~A | ~B) & (~A | B)

endmodule
