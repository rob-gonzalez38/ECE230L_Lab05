module circuit_b(
    // Declare inputs
    // Declare Y output
);

    // Enter logic equation here
    (~C & ~D) | (A & B) | (B & C & ~D)

endmodule
